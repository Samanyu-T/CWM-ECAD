//////////////////////////////////////////////////////////////////////////////////
// Test bench for Exercise #8  - Simple End-to-End Design
// Student Name:
// Date: 
//
// Description: A testbench module to test Ex8
// You need to write the whole file
//////////////////////////////////////////////////////////////////////////////////

//I don't have enough time to fully write this so:
//Make registers to store the inputs to top.v, i.e reg temperature_0 = 1'b0 and so on 
//Not sure on how to input the clock signals 
//Once this is intialise simply use the same test criterion as in Excercise 5
//So send 1 set of data and check if the output is reasonable.
